`timescale 1ns / 1ps
`default_nettype none
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/20/2019 04:26:22 PM
// Design Name: 
// Module Name: phywhisperer_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module tb_pw();
   
    parameter pUSB_CLOCK_PERIOD = 10;
    parameter pFE_CLOCK_PERIOD = 16;
    // TODO: generate a few testcases wih various ranges of delays, to more easily stress and hit corner cases
    parameter pMIN_FE_DELAY = 0;
    parameter pMAX_FE_DELAY = 7;
    parameter pDELAY_MODE = 0;
    parameter pVERBOSE = 1;
    parameter pNUM_EVENTS = 20;
    parameter pSEED = 1;

   // FIFO bitfields: (TODO: pull in from external file)
   `define FE_FIFO_CMD_DATA 2'b00
   `define FE_FIFO_CMD_STAT 2'b01
   `define FE_FIFO_CMD_TIME 2'b10

   `define FE_FIFO_CMD_START 16
   `define FE_FIFO_CMD_BIT_LEN 2

   `define FE_FIFO_TIME_START 0
   `define FE_FIFO_SHORTTIME_LEN 3
   `define FE_FIFO_FULLTIME_LEN 16

   `define FE_FIFO_RXACTIVE_BIT 3
   `define FE_FIFO_RXERROR_BIT 4
   `define FE_FIFO_SESSVLD_BIT 5
   `define FE_FIFO_SESSEND_BIT 6
   `define FE_FIFO_VBUSVLD_BIT 7

   `define FE_FIFO_DATA_START 8
   `define FE_FIFO_DATA_LEN 8


    reg           usb_clk;
    wire [7:0]    USB_Data;
    reg  [7:0]    USB_wdata;
    reg  [7:0]    USB_Addr;
    reg           USB_nRD;
    reg           USB_nWE;
    reg           USB_nCS;
    wire          USB_SPARE0;
    reg           USB_SPARE1;

    /* FRONT END CONNECTIONS */
    reg  fe_clk;
    reg  fe_txrdy;
    reg  fe_rxactive;
    reg  fe_id_dig;
    reg  fe_linestate0;
    reg  fe_linestate1;
    reg  fe_hostdisc;
    reg  fe_sessend;
    wire [7:0] fe_data;
    reg  [7:0] fe_wdata;
    reg  fe_rxvalid;
    reg  fe_sessvld;
    reg  fe_rxerror;
    reg  fe_vbusvld;

    /* 20-PIN USER HEADER CONNECTOR */
    reg  [7:0] userio_d;
    reg  userio_clk;
    reg  [23:0] read_data;
    reg  [7:0] data;
    reg  [1:0] command;
    reg  [`FE_FIFO_FULLTIME_LEN-1:0] timestamp;

    /* 20-PIN CHIPWHISPERER CONNECTOR */
    wire cw_clk;
    wire cw_trig;

    reg  reset;
    int  seed;


    //TODO: provide input seed, so user running testbench can choose to change it or repeat it

   initial begin
      seed = pSEED;
      $display("Running with pSEED=%0d", pSEED);
      $urandom(seed);
      $dumpfile("tb.fst");
      $dumpvars(0, tb_pw);
      usb_clk = 1'b1;
      fe_clk = 1'b1;
      reset = 1'b0;

      USB_wdata = 0;
      USB_Addr = 0;
      USB_nRD = 1;
      USB_nWE = 1;
      USB_nCS = 1;
      USB_SPARE1 = 1;

      fe_txrdy = 0;
      fe_rxactive = 0;
      fe_id_dig = 0;
      fe_linestate0 = 0;
      fe_linestate1 = 0;
      fe_hostdisc = 0;
      fe_sessend = 0;
      fe_wdata = 0;
      fe_rxvalid = 0;
      fe_sessvld = 0;
      fe_rxerror = 0;
      fe_vbusvld = 0;

      //userio_d = 0;
      //userio_clk = 0;

      #(pUSB_CLOCK_PERIOD*2) reset = 1;
      #(pUSB_CLOCK_PERIOD*2) reset = 0;

      /*
      repeat(10) @(posedge usb_clk);
      write_1byte(0, 8'ha3);
      repeat(10) @(posedge usb_clk);
      read_1byte(0, read_data);
      $display("Got %h", read_data);
      */

      //#(pFE_CLOCK_PERIOD*100) $finish;
   end

   int i,j;
   int errors;
   int time_counter;
   reg [7:0] fe_bytes [0:2047];
   reg [15:0] fe_times [0:2047];

   // FE feeding thread:
   initial begin
      errors = 0;
      #(pFE_CLOCK_PERIOD*100);
      write_1byte(2, 8'h01); // enable timestamps
      write_1byte(3, 8'h01); // enable capture
      fe_times[0] = 0; // by definition

      if (pVERBOSE) begin
         $display("------------------------------|-------------------------------");
         $display("FE testbench sending:         | PhyWhisperer DUT receiving:");
         $display("------------------------------|-------------------------------");
      end

      @(posedge fe_clk);
      for (i = 0; i < pNUM_EVENTS; i = i + 1) begin
         fe_bytes[i] = $urandom;
         get_delay(fe_times[i+1]);
         send_fe_data(fe_bytes[i], fe_times[i+1]);
         if (pVERBOSE)
            $display("data=%h, delay=%0d", fe_bytes[i], fe_times[i+1]);
      end
      fe_rxvalid = 1'b0;
      #(pFE_CLOCK_PERIOD*1000);
      if (j == pNUM_EVENTS)
         $display("Read all %0d DATA packets", j);
      else begin
         $display("*** ONLY READ %0d of %0d DATA packets.", j, pNUM_EVENTS);
         errors += 1;
      end
      if (errors)
         $display("SIMULATION FAILED (%0d errors).", errors);
      else
         $display("Simulation passed!");
      $finish;
   end


   // FIFO read thread:
   initial begin
      j = 0;
      time_counter = 0;
      while (1) begin
         wait (U_dut.U_reg_pw.sniff_fifo_empty == 1'b0);
         read_lots_bytes(1);
         read_next_byte(read_data[7:0]);
         read_next_byte(read_data[15:8]);
         read_next_byte(read_data[23:16]);
         command = read_data[`FE_FIFO_CMD_START +: `FE_FIFO_CMD_BIT_LEN];

         if (command == `FE_FIFO_CMD_DATA) begin
            data = read_data[`FE_FIFO_DATA_START +: `FE_FIFO_DATA_LEN];
            timestamp = read_data[`FE_FIFO_TIME_START +: `FE_FIFO_SHORTTIME_LEN];
            time_counter = time_counter + timestamp;
            if ( (data == fe_bytes[j]) && (time_counter == fe_times[j]) ) begin
               if (pVERBOSE)
                  $display("\t\t\t\tdata=%h, time=%0d, total time=%0d", data, timestamp, time_counter);
            end
            else begin
               errors += 1;
               if (data == fe_bytes[j])
                  $display("\t\t\t\t*** MISMATCH on FIFO read #%0d at time %0t: got good data (%h), bad time: expected %0d, got %0d (DATA time=%0d)", j, $time, data, fe_times[j], time_counter, timestamp);
               else if (time_counter == fe_times[j])
                  $display("\t\t\t\t*** MISMATCH on FIFO read #%0d at time %0t: got good timestamp (%0d), bad data: got %h, expected %h", j, $time, timestamp, data, fe_bytes[j]);
               else
                  $display("\t\t\t\t*** MISMATCH on FIFO read #%0d at time %0t: bad data (got %h, expected %h) and bad time (got %0d, expecte %0d)", j, $time, data, fe_bytes[j], time_counter, fe_times[j]);
            end
            j = j + 1;
            time_counter = 0;
         end

         else if (command == `FE_FIFO_CMD_STAT) begin
            $display("\t\t\t\t*** ERROR: STAT command not supported yet!");
         end

         else if (command == `FE_FIFO_CMD_TIME) begin
            timestamp = read_data[`FE_FIFO_TIME_START +: `FE_FIFO_FULLTIME_LEN];
            time_counter = time_counter + timestamp;
            if (pVERBOSE)
               $display("\t\t\t\ttime=%0d", timestamp);
         end

         else begin
            errors += 1;
            $display("\t\t\t\t*** ERROR: Unknown command!");
         end

      end
   end


   assign USB_Data = USB_nWE? 8'bz : USB_wdata;
   assign fe_data = fe_wdata;
   assign USB_SPARE0 = reset;

   task write_1byte;
      input [7:0] address;
      input [7:0] data;
      @(posedge usb_clk);
      USB_SPARE1 = 0;
      USB_Addr = address;
      @(posedge usb_clk);
      USB_SPARE1 = 1;
      repeat(4) @(posedge usb_clk);
      USB_wdata = data;
      USB_nWE = 0;
      @(posedge usb_clk);
      USB_nWE = 1;
      USB_nCS = 0;
      @(posedge usb_clk);
      USB_nCS = 1;
   endtask


   task read_1byte;
      input [7:0] address;
      output [7:0] data;
      @(posedge usb_clk);
      USB_SPARE1 = 0;
      USB_Addr = address;
      @(posedge usb_clk);
      USB_SPARE1 = 1;
      repeat(4) @(posedge usb_clk);
      USB_nRD = 0;
      USB_nCS = 0;
      @(posedge usb_clk);
      USB_nCS = 1;
      //data = USB_Data;
      @(posedge usb_clk);
      #1 data = USB_Data;
      @(posedge usb_clk);
      USB_nRD = 1;
   endtask

   task read_lots_bytes;
      input [7:0] address;
      @(posedge usb_clk);
      USB_SPARE1 = 0;
      USB_Addr = address;
      @(posedge usb_clk);
      USB_SPARE1 = 1;
      repeat(4) @(posedge usb_clk);
   endtask

   task read_next_byte;
      output [7:0] data;
      USB_nRD = 0;
      USB_nCS = 0;
      @(posedge usb_clk);
      USB_nCS = 1;
      @(posedge usb_clk);
      #1 data = USB_Data;
      @(posedge usb_clk);
      USB_nRD = 1;
      @(posedge usb_clk);
   endtask


   task send_fe_data;
      input [7:0] data;
      input [15:0] delay;
      fe_rxvalid = 1;
      fe_wdata = data;
      @(posedge fe_clk);
      if (delay > 0) begin
         fe_rxvalid = 0;
         fe_wdata = 0;
      end
      repeat (delay) @(posedge fe_clk);
   endtask


   task get_delay;
      output [15:0] delay;
      if (pDELAY_MODE == 0)
         delay = $urandom_range(pMIN_FE_DELAY, pMAX_FE_DELAY);
      else if (pDELAY_MODE == 1) begin
         delay = $urandom_range(0, 1);
         if (delay == 1) delay = $urandom_range(pMIN_FE_DELAY, pMAX_FE_DELAY);
         else delay = 0;
      end
   endtask



   always #(pUSB_CLOCK_PERIOD/2) usb_clk = !usb_clk;
   always #(pFE_CLOCK_PERIOD/2) fe_clk = !fe_clk;

   // TODO: repeat this for all DUT inputs
   wire #1 fe_id_dig_out      = fe_id_dig;
   wire #1 fe_txrdy_out       = fe_txrdy;
   wire #1 fe_rxactive_out    = fe_rxactive;
   wire #1 fe_linestate0_out  = fe_linestate0;
   wire #1 fe_linestate1_out  = fe_linestate1;
   wire #1 fe_hostdisc_out    = fe_hostdisc;
   wire #1 fe_sessend_out     = fe_sessend;
   wire [7:0] #1 fe_data_out  = fe_data;
   wire #1 fe_rxvalid_out     = fe_rxvalid;
   wire #1 fe_sessvld_out     = fe_sessvld;
   wire #1 fe_rxerror_out     = fe_rxerror;
   wire #1 fe_vbusvld_out     = fe_vbusvld;

phywhisperer_top U_dut (
    /* USB CHIP CONNECTIONS */
    .usb_clk            (usb_clk    ),
    .USB_Data           (USB_Data   ),
    .USB_Addr           (USB_Addr   ),
    .USB_nRD            (USB_nRD    ),
    .USB_nWE            (USB_nWE    ),
    .USB_nCS            (USB_nCS    ),
    .USB_SPARE0         (USB_SPARE0 ),
    .USB_SPARE1         (USB_SPARE1 ),

    /* FRONT END CONNECTIONS */
    .fe_xcvrsel0        (), // unused
    .fe_xcvrsel1        (), // unused
    .fe_termsel         (), // unused
    .fe_suspendn        (), // unused
    .fe_txvalid         (), // unused
    .fe_reset           (), // unused
    .fe_chrgvbus        (), // unused
    .fe_opmode0         (), // unused
    .fe_opmode1         (), // unused
    .fe_idpullup        (), // unused
    .fe_dischrgvbus     (), // unused
    .fe_dppd            (), // unused
    .fe_dmpd            (), // unused
    .fe_id_dig          (fe_id_dig_out     ),
    .fe_txrdy           (fe_txrdy_out      ),
    .fe_rxactive        (fe_rxactive_out   ),
    .fe_linestate0      (fe_linestate0_out ),
    .fe_linestate1      (fe_linestate1_out ),
    .fe_hostdisc        (fe_hostdisc_out   ),
    .fe_sessend         (fe_sessend_out    ),
    .fe_clk             (fe_clk            ),
    .fe_data            (fe_data_out       ),
    .fe_rxvalid         (fe_rxvalid_out    ),
    .fe_sessvld         (fe_sessvld_out    ),
    .fe_rxerror         (fe_rxerror_out    ),
    .fe_vbusvld         (fe_vbusvld_out    ),

    /* 20-PIN USER HEADER CONNECTOR */
    .userio_d           (userio_d),
    .userio_clk         (userio_clk),

    /* 20-PIN CHIPWHISPERER CONNECTOR */
    .cw_clk             (cw_clk),
    .cw_trig            (cw_trig)
    );

endmodule
`default_nettype wire

